------------------------------------------------------------------------------
-- Name : 
-- Last Update : 
-- Tested : 
--
-- Desc : Bla bli blo
------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

--library work;
--use work.pkg_parameters.all;


entity <name> is
    Port ( 

    ); 
end <name> ;


architecture rtl of <name>  is

    ---------------
    -- CONSTANTS --
    ---------------

    -----------
    -- TYPES --
    -----------

    -------------
    -- SIGNALS --
    -------------

begin

    -- Input (Optional)


    -- Output

end architecture;